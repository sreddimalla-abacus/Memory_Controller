class mem_mon;
  task run();
    $display("mem_mon::run");
  endtask
endclass