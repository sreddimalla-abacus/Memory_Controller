program mc_tb();
  mc_env env;
  initial begin
    env = new();
    env.run();
    
  end
endprogram
