class wb_mon;
  task run();
    $display("wb_mon::run");
  endtask
endclass