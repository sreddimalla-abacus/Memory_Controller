class mc_ref;
  task run();
    $display("mc_ref::run");
  endtask
endclass