class mc_ckr;
  task run();
    $display("mc_ckr::run");
  endtask
endclass