class wb_cov;
  task run();
    $display("wb_cov::run");
  endtask
endclass